
module imm_gen #(parameter  mode=32 )(
    input [mode-1 : 0]instruction,
    output [mode-1 : 0]imm
);

always_comb begin
    

    
    
end



endmodule
